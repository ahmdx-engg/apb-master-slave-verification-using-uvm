package tx_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  // List components in dependency order
  // `include "agent_config.sv"
  `include "tx_item.sv"
  `include "first_sequence.sv"
  `include "sequencer.sv"
  `include "monitor.sv"
  `include "driver.sv"
  `include "agent.sv"
  `include "scoreboard.sv"
  // `include "evaluator.sv"
  `include "env.sv"
  `include "test.sv"
endpackage